-- Author(s):     Nuttanon Pongpunlux 6538050421
--                Siraphop Wannasanmethar 6538213421
--                Supadet Udomgewganchana 6538205421
--
-- Date:          10 May 2025
--
-- Description:
--    Logic Design (2147307) Final Project
--    Full Adder component implemented with multiple architectures:
--    1. Logic equations
--    2. Half adder-based
--    3. Multiplexer-based
--    4. Numeric-based (for synthesis readability)

-- Standard library inclusions
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.std_logic_misc.ALL;
USE IEEE.vital_timing.ALL;  -- Provides timing delay definitions

-- Entity for full adder with timing delay parameters
ENTITY full_adder IS
    GENERIC (
        -- Timing parameters (in nanoseconds)
        tpd_x_s       : TIME := 1 ns;  -- Delay from input x to output s
        tpd_y_s       : TIME := 1 ns;  -- Delay from input y to output s
        tpd_cin_s     : TIME := 1 ns;  -- Delay from carry-in to sum
        tpd_x_cout    : TIME := 1 ns;  -- Delay from x to carry-out
        tpd_y_cout    : TIME := 1 ns;  -- Delay from y to carry-out
        tpd_cin_cout  : TIME := 1 ns   -- Delay from carry-in to carry-out
    );
    PORT (
        Cin   : IN  STD_LOGIC;  -- Carry-in input
        x     : IN  STD_LOGIC;  -- Operand 1
        y     : IN  STD_LOGIC;  -- Operand 2
        s     : OUT STD_LOGIC;  -- Sum output
        Cout  : OUT STD_LOGIC   -- Carry-out output
    );

    -- Design documentation:
    -- A full adder adds three bits: x, y, and Cin.
    -- Produces: sum (s) and carry-out (Cout)
    -- Truth table:
    --   x y Cin | s Cout
    --   0 0 0   | 0  0
    --   0 0 1   | 1  0
    --   0 1 0   | 1  0
    --   0 1 1   | 0  1
    --   1 0 0   | 1  0
    --   1 0 1   | 0  1
    --   1 1 0   | 0  1
    --   1 1 1   | 1  1
END ENTITY full_adder;

--===========================================================
-- Architecture 1: Logic equations
--===========================================================
ARCHITECTURE LogicFunc OF full_adder IS
BEGIN
    -- Standard equation for sum: XOR all three inputs
    s    <= x XOR y XOR Cin AFTER tpd_x_s;

    -- Carry-out is generated by majority function of inputs
    Cout <= (x AND y) OR (Cin AND x) OR (Cin AND y) AFTER tpd_x_cout;
END ARCHITECTURE LogicFunc;

--===========================================================
-- Architecture 2: Using two half adders
--===========================================================
ARCHITECTURE HalfAdders OF full_adder IS
    SIGNAL sum1, carry1, carry2 : STD_LOGIC;  -- Intermediate signals
BEGIN
    -- First half adder: x + y
    sum1   <= x XOR y AFTER tpd_x_s;
    carry1 <= x AND y AFTER tpd_x_cout;

    -- Second half adder: sum1 + Cin
    s      <= sum1 XOR Cin AFTER tpd_cin_s;
    carry2 <= sum1 AND Cin AFTER tpd_cin_cout;

    -- Final carry is OR of both half adder carries
    Cout   <= carry1 OR carry2 AFTER 0.5 ns;
END ARCHITECTURE HalfAdders;

--===========================================================
-- Architecture 3: Optimized with multiplexer logic
--===========================================================
ARCHITECTURE Optimized OF full_adder IS
BEGIN
    -- XOR remains for sum
    s <= x XOR y XOR Cin AFTER tpd_x_s;

    -- Optimized carry: if x = y, Cout = x; else Cout = Cin
    Cout <= x WHEN (x = y) ELSE Cin AFTER tpd_x_cout;
END ARCHITECTURE Optimized;

--===========================================================
-- Architecture 4: Using integer-based logic (good for synthesis)
--===========================================================
ARCHITECTURE Numeric OF full_adder IS
    SIGNAL temp_sum : INTEGER RANGE 0 TO 3;  -- Sum of 3 input bits
BEGIN
    -- Integer-based input encoding
    temp_sum <= 0 WHEN x = '0' AND y = '0' AND Cin = '0' ELSE
                1 WHEN (x = '1' AND y = '0' AND Cin = '0') OR
                      (x = '0' AND y = '1' AND Cin = '0') OR
                      (x = '0' AND y = '0' AND Cin = '1') ELSE
                2 WHEN (x = '1' AND y = '1' AND Cin = '0') OR
                      (x = '1' AND y = '0' AND Cin = '1') OR
                      (x = '0' AND y = '1' AND Cin = '1') ELSE
                3;

    -- Output based on integer sum
    s    <= '1' WHEN (temp_sum = 1) OR (temp_sum = 3) ELSE '0' AFTER tpd_x_s;
    Cout <= '1' WHEN (temp_sum >= 2) ELSE '0' AFTER tpd_x_cout;
END ARCHITECTURE Numeric;
